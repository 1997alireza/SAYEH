library IEEE;
use IEEE.std_logic_1164.all;

entity CU is

end entity;

architecture CU_ARCH of CU is 
begin
  
end architecture;




